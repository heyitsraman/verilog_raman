// Hello World Example
module hello_world();
    initial begin
      $display("\n\t Hello World! This is Revti Raman. \n");
    end

endmodule